
/*
 *  tISRWithInterruptRequest �� celltype �L�q
 */
import("Temp.cdl");

/* �R�[���o�b�N���[�`���̎��ʔԍ� */
const uint_t SIO_RDY_SND = 1;		/* ���M�\�R�[���o�b�N */
const uint_t SIO_RDY_RCV = 2;		/* ��M�ʒm�R�[���o�b�N */

celltype tSIOPortSkyeyeMain {
	entry sSIOPort	eSIOPort;
	call siSIOCBR	ciSIOCBR;

	entry sRoutineBody eInitialize; /* ���������� */
	entry sRoutineBody eTerminate;  /* �I������ */

	entry siHandlerBody eiISR;/* �����݃T�[�r�X���[�`�� */
	
	attr {
		/*Skyeye�p�̃A�h���X*/
		uint32_t  uartBase;
	};
	var {
		/*
		 * skyeye�p
		 */
		bool_t	openFlag;			/* �I�[�v���ς݃t���O */
		bool_t	receiveFlag;			/* ��M�����o�b�t�@�L���t���O */
		char_t	receiveBuffer;			/* ��M�����o�b�t�@ */
		bool_t	receiveReady;			/* ��M�ʒm�R�[���o�b�N���t���O */
		/* SkyEye�̏ꍇ�͑��M�͏�ɂł���̂ŁA���M�����o�b�t�@�͕K�v�Ȃ� */
     	bool_t	sendReady;			/* ���M�ʒm�R�[���o�b�N���t���O */
	};
	FACTORY {
		write("$ct$_factory.h", "#include \"at91skyeye.h\"");
	};
};

[active]
composite tSIOPortSkyeye {
	entry sSIOPort	eSIOPort;
	call siSIOCBR	ciSIOCBR;

	attr {
		/*Skyeye�p�̃A�h���X*/
		//uint32_t* uartBase = C_EXP("(USART0_BASE)");
		uint32_t uartBase = 0xFFFD0000;
	};

	cell tSIOPortSkyeyeMain SIOPortMain {
		ciSIOCBR => composite.ciSIOCBR;
		uartBase = composite.uartBase;
	};
	/*
	 *  �Ȉ�SIO�h���C�o�̏������������[�`��
	 */
	cell tInitializeRoutine InitializeSIO{
		cInitializeRoutineBody = SIOPortMain.eInitialize;
	};
	/*
	 *  �Ȉ�SIO�h���C�o�̏I���������[�`��
	 */
	cell tTerminateRoutine TerminateSIO{
		cTerminateRoutineBody = SIOPortMain.eTerminate;
	};
	cell tISRWithInterruptRequest SIOPortSkyeyeISR{
		ciISRBody =  SIOPortMain.eiISR;
		interruptNumber   =  2;
		interruptPriority = -2;
	};
	composite.eSIOPort => SIOPortMain.eSIOPort;
};
	
