/*
 * 
 */
[singleton]
celltype tPutLogSkyeye {
	entry sPutLog	ePutLog;
	call  sSIOPort  cSIOPort;
};
