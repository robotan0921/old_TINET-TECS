 /*
  * ��ˑ����ɒ񋟂���֐�
  */
signature sSIOPort {
 	void	open(void);
	void	close(void);
	bool_t	putChar([in] char_t c);
	int_t	getChar(void);
	void	enableCBR([in] uint_t cbrtn);
	void	disableCBR([in] uint_t cbrtn);
};
/*
 * ��ˑ����ւ̃R�[���o�b�N
 */
signature siSIOCBR {
	void	readySend(void);
	void	readyReceive(void);
};

/* �R�[���o�b�N���[�`���̎��ʔԍ� */
const uint_t SIO_RDY_SND = 1;		/* ���M�\�R�[���o�b�N */
const uint_t SIO_RDY_RCV = 2;		/* ��M�ʒm�R�[���o�b�N */

celltype tSIOPortSkyeyeMain {
	entry sSIOPort	eSIOPort;
	call siSIOCBR	ciSIOCBR;

	entry sInitializeRoutineBody eInitialize; /* ���������� */
	entry sTerminateRoutineBody eTerminate;   /* �I������ */

	entry siHandlerBody eiISR;/* �����݃T�[�r�X���[�`�� */
	
	attr {
		/*Skyeye�p�̃A�h���X*/
		uint32_t  uartBase;
	};
	var {
		/*
		 * skyeye�p
		 */
		bool_t	openFlag;			/* �I�[�v���ς݃t���O */
		bool_t	receiveFlag;			/* ��M�����o�b�t�@�L���t���O */
		char_t	receiveBuffer;			/* ��M�����o�b�t�@ */
		bool_t	receiveReady;			/* ��M�ʒm�R�[���o�b�N���t���O */
		/* SkyEye�̏ꍇ�͑��M�͏�ɂł���̂ŁA���M�����o�b�t�@�͕K�v�Ȃ� */
     	bool_t	sendReady;			/* ���M�ʒm�R�[���o�b�N���t���O */
	};
	FACTORY {
		write("$ct$_factory.h", "#include \"at91skyeye.h\"");
	};
};

[active]
composite tSIOPortSkyeye {
	entry sSIOPort	eSIOPort;
	call siSIOCBR	ciSIOCBR;

	attr {
		/*Skyeye�p�̃A�h���X*/
		//uint32_t* uartBase = C_EXP("(USART0_BASE)");
		uint32_t uartBase = 0xFFFD0000;
	};

	cell tSIOPortSkyeyeMain SIOPortMain {
		ciSIOCBR => composite.ciSIOCBR;
		uartBase = composite.uartBase;
	};
	/*
	 *  �Ȉ�SIO�h���C�o�̏������������[�`��
	 */
	cell tInitializeRoutine InitializeSIO{
		cInitializeRoutine = SIOPortMain.eInitialize;
	};
	/*
	 *  �Ȉ�SIO�h���C�o�̏I���������[�`��
	 */
	cell tTerminateRoutine TerminateSIO{
		cTerminateRoutine = SIOPortMain.eTerminate;
	};
	cell tISRWithConfigInterrupt SIOPortSkyeyeISR{
		ciBody =  SIOPortMain.eiISR;
		interruptNumber   =  2;
		interruptPriority = -2;
	};
	composite.eSIOPort => SIOPortMain.eSIOPort;
};
	