/*     �C�[�T�l�b�g�o�̓^�X�N
          ID�FETHER_OUTPUT_TASK
          �D��x�F5
          ������ԁFTA_HLNG
          �ďo���֐��Fehter_output_task(net/ethernet.c)
          �X�^�b�N�T�C�Y�F1024
     �C�[�T�l�b�g���̓^�X�N
          ID�FETHER_INPUT_TASK
          �D��x�F5
          ������ԁFTA_HLNG
          �ďo���֐��Fehter_input_task(net/ethernet.c)
          �X�^�b�N�T�C�Y�F1024         
*/





signature sArpInput{
    void arpInitialize(void);
    void arpInput([send(sNetworkAlloc),size_is(size)] int8_t *inputp,[in]int32_t size,[in,size_is(6)]const uint8_t *macaddress);
};

signature sIPv4Input {
    void IPv4Input([send(sNetworkAlloc),size_is(size)] int8_t *inputp,[in]int32_t size);
};


celltype tEthernetInputTaskBody {

    call sSemaphore cSemaphoreReceive;
    call sNicDriver cNicDriver;
    
    [optional]call sTask cTaskEthernetOutput;
    call sTask cTaskNetworkTimer;

    [optional]call sArpInput cArpInput;
    [optional]call sIPv4Input cIPv4Input;

    entry sTaskBody eBody;
};






signature sEthernetRawOutput{
    ER ethernetRawOutput([send(sNetworkAlloc),size_is(size)]int8_t *outputp,[in]int32_t size,[in]TMO tmout);
};

signature sArpOutput{
    ER arpResolve([send(sNetworkAlloc),size_is(size)] int8_t *outputp,[in]int32_t size,[in]T_IN4_ADDR dstaddr,[in,size_is(6)]const uint8_t *macaddress,[in]TMO tmout);
};

signature sEthernetOutput{
    ER ethernetOutput([send(sNetworkAlloc),size_is(size)] int8_t *outputp,[in]int32_t size,[in]T_IN4_ADDR dstaddr,[in]TMO tmout);
};
    
celltype tEthernetOutput {
    call sEthernetRawOutput cRawOutput;
    call sNicDriver cNicDriver;
    [optional]call sArpOutput cArpOutput;

    entry sEthernetOutput eEthernetOutput;
};


celltype tEthernetOutputTaskBody {

    require tKernel.eKernel;

    call sSemaphore cSemaphoreSend;
    call sDataqueue cDataqueue;
    call sNicDriver cNicDriver;

    [optional]call sSemaphore cSemTcppost;

    entry sEthernetRawOutput eRawOutput;
    entry sTaskBody eBody;
};

/*�R���|�W�b�g�����̃Z���h���V�[�u���g���Ȃ�
[active]
composite tEthernetOutputComposite{

    attr{
        uint_t countQueue;
        PRI taskPriority;
        SIZE taskSize;
    };

    call sNicDriver cNicDriver;
    call sSemaphore cSemaphoreSend;
    [optional]call sArpOutput cArpOutput;

    entry sTask eEthernetOutputTask;
    entry sEthernetRawOutput eRawOutput;
    entry sEthernetOutput eEthernetOutput;
    

    cell tDataqueue Dataqueue{
        attribute = C_EXP("TA_NULL");
        count = composite.countQueue;
        pdqmb = C_EXP("NULL");
    };

    [allocator(eRawOutput.ethernetRawOutput.output=NetworkBuffer.eNetworkAlloc)]
    cell tEthernetOutputTaskBody EthernetOutputTaskBody{
        cNicDriver => composite.cNicDriver;
        cSemaphoreSend =>composite.cSemaphoreSend;
        cDataqueue = Dataqueue.eDataqueue;
    };
    
    cell tTask Task{
        cBody = EthernetOutputTaskBody.eBody;

        taskAttribute = C_EXP("TA_NULL");
        priority = taskPriority;
        stackSize = taskSize;
    };

    cell tEthernetOutput EthernerOutput{
        cRawOutput = EthernetOutputTaskBody.eRawOutput;
        cArpOutput => composite.cArpOutput;
        cNicDriver => composite.cNicDriver;
    };

    composite.eEthernetOutputTask => Task.eTask;
    composite.eRawOutput => EthernetOutputTaskBody.eRawOutput;
    composite.eEthernetOutput => EthernerOutput.eEthernetOutput;
};
  */