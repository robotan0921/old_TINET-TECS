
signature sTINET{
    uint32_t netRand(void);
    void netSrand([in]uint32_t speed);
};
    

[singleton]
celltype tTINET{
    var{
        uint32_t next = 1;
    };

    entry sTINET eTINET;
};


//�l�b�g���[�N�p�������A���P�[�^�̒�`�ƃZ����
import ("tBuffer.cdl");

//�e�w���Ƃ̃}�N����`
import_C ("tecsinet.h");
import_C ("Ethernet_define.h");
import_C("ipv4_define.h");
import_C("ipv6_define.h");
import_C("udp_define.h");
import_C("tcp_define.h");


//�l�b�g���[�N�^�C�}�R���|�[�l���g�̒�`
import ("tNetworkTimer.cdl");



//Lan9221�p�f�o�h���R���|�[�l���g�̒�`
import ("tLan9221.cdl");

//Ethernet���C���p�̃R���|�[�l���g��`����
import ("tEthernet.cdl");

//IPv4���C���p�̃R���|�[�l���g��`����
import ("tIPv4.cdl");

//IPv6���C���p�̃R���|�[�l���g��`����
import ("tIPv6.cdl");

//UDP���C���p�̃R���|�[�l���g��`����
import ("tUDP.cdl");

//TCP���C���p�̃R���|�[�l���g��`����
import ("tTCP.cdl");
