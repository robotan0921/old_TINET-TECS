//************************************************

//            ��`

//************************************************

//�ڑ����Ă���^�C�}�[�֐�(���߂ł�OK���j
const uint32_t NUM_NETWORKTIMER=5;

//�^�C�}�̋O������
const uint32_t NET_TIMER_CYCLE=100;

//�^�C�}�^�X�N�̗D��x
const int32_t NET_TIMER_PRIORITY=3;


//************************************************

//            �Z���^�C�v�錾

//************************************************


[singleton]
celltype tNetworkTimer{
    /*attr{
        [size_is(NUM_NETWORKTIMER)]int32_t *timeoutTemp;
    };*/
    var {
        [size_is(NUM_NETWORKTIMER)]int32_t *timeout = {-1,-1,-1,-1};
    };

    [optional]call sCallTimerFunction cCallTimerFunction[NUM_NETWORKTIMER];

    [optional]call sTask cTCPTask;

    call sSemaphore cSemaphoreNetworkTimer;
    call siSemaphore ciSemaphoreNetworkTimer;
    call sSemaphore cSemaphoreCalloutLock;

    entry sNetworkTimer eNetworkTimer[NUM_NETWORKTIMER];


    entry sTaskBody eBody;
    entry siHandlerBody eiBody;
};


//************************************************

//            �g�ݏグ�錾

//************************************************


cell tNetworkTimer NetworkTimer;


cell tCyclicHandler NetTimerHandler{
    ciBody = NetworkTimer.eiBody;
    
    attribute = C_EXP("TA_ACT");
    cyclicTime = NET_TIMER_CYCLE;
    cyclicPhase = 1;
};

cell tTask NetTimerTask{
    cBody = NetworkTimer.eBody;

    taskAttribute = C_EXP("TA_NULL");
    priority = NET_TIMER_PRIORITY;
    stackSize = 1024;
};

cell tSemaphore SemaphoreNetworkTimer{
    attribute = C_EXP("TA_TPRI");
    count = 0;
    max = NUM_NETWORKTIMER;
};

cell tSemaphore SemaphoreCalloutLock{
    attribute = C_EXP("TA_TPRI");
    count = 1;
    max = 1;
};